library ieee;
use ieee.std_logic_1164.all;

entity Aktivno_stanje is
	port(
		enable: in std_logic
	);
end Aktivno_stanje;

architecture Beh of Aktivno_stanje is


begin

end Beh;