library verilog;
use verilog.vl_types.all;
entity Ploca_B_vlg_vec_tst is
end Ploca_B_vlg_vec_tst;
